module clockdivider(
	input logic reset,
	output logic clk,
	output logic [10:0] counter
);
	logic int_osc;

	// Internal high-speed oscillator
	HSOSC hf_osc (.CLKHFPU(1'b1), .CLKHFEN(1'b1), .CLKHF(int_osc));
	
	// Simple clock divider
	always_ff @(posedge int_osc) begin
		if (reset==0) 	counter = 0;
		else 		counter = counter + 1;
		end
	assign clk = counter[10];
endmodule